<svg width="297mm" height="420mm" viewBox="0 0 1122 1587" xmlns="http://www.w3.org/2000/svg">
  <defs>
    <!-- Gradients for cosmic background -->
    <radialGradient id="cosmicBg" cx="50%" cy="30%" r="70%">
      <stop offset="0%" style="stop-color:#1a0033;stop-opacity:0.8"/>
      <stop offset="30%" style="stop-color:#2d1b69;stop-opacity:0.7"/>
      <stop offset="70%" style="stop-color:#0f0520;stop-opacity:0.8"/>
      <stop offset="100%" style="stop-color:#000000;stop-opacity:0.9"/>
    </radialGradient>
    
    <!-- Planet glows -->
    <filter id="glow" x="-50%" y="-50%" width="200%" height="200%">
      <feGaussianBlur stdDeviation="8" result="coloredBlur"/>
      <feMerge> 
        <feMergeNode in="coloredBlur"/>
        <feMergeNode in="SourceGraphic"/>
      </feMerge>
    </filter>
    
    <filter id="strongGlow" x="-100%" y="-100%" width="300%" height="300%">
      <feGaussianBlur stdDeviation="15" result="coloredBlur"/>
      <feMerge> 
        <feMergeNode in="coloredBlur"/>
        <feMergeNode in="SourceGraphic"/>
      </feMerge>
    </filter>
    
    <!-- Spaceship thruster animation -->
    <radialGradient id="thruster" cx="50%" cy="50%" r="50%">
      <stop offset="0%" style="stop-color:#00ffff;stop-opacity:1">
        <animate attributeName="stop-opacity" values="1;0.3;1" dur="0.5s" repeatCount="indefinite"/>
      </stop>
      <stop offset="50%" style="stop-color:#0066ff;stop-opacity:0.8">
        <animate attributeName="stop-opacity" values="0.8;0.2;0.8" dur="0.5s" repeatCount="indefinite"/>
      </stop>
      <stop offset="100%" style="stop-color:#003366;stop-opacity:0"/>
    </radialGradient>
    
    <!-- Path gradient -->
    <linearGradient id="pathGrad" x1="0%" y1="0%" x2="100%" y2="100%">
      <stop offset="0%" style="stop-color:#00ffff;stop-opacity:0.8"/>
      <stop offset="50%" style="stop-color:#ff6600;stop-opacity:0.6"/>
      <stop offset="100%" style="stop-color:#ff0066;stop-opacity:0.8"/>
    </linearGradient>
    
    <!-- Star twinkle animation -->
    <animate id="twinkle" attributeName="opacity" values="0.3;1;0.3" dur="2s" repeatCount="indefinite"/>
  </defs>
  
  <!-- Cosmic background -->
  <rect width="100%" height="100%" fill="url(#cosmicBg)"/>
  
  <!-- Stars -->
  <circle cx="150" cy="200" r="1.5" fill="#ffffff" opacity="0.8">
    <use href="#twinkle"/>
  </circle>
  <circle cx="300" cy="150" r="1" fill="#ffff99" opacity="0.6">
    <animate attributeName="opacity" values="0.6;1;0.6" dur="3s" repeatCount="indefinite"/>
  </circle>
  <circle cx="450" cy="180" r="1.2" fill="#ffffff" opacity="0.7">
    <use href="#twinkle"/>
  </circle>
  <circle cx="600" cy="120" r="1" fill="#99ccff" opacity="0.5">
    <animate attributeName="opacity" values="0.5;0.9;0.5" dur="2.5s" repeatCount="indefinite"/>
  </circle>
  <circle cx="750" cy="200" r="1.3" fill="#ffffff" opacity="0.8">
    <use href="#twinkle"/>
  </circle>
  <circle cx="900" cy="160" r="1" fill="#ffccff" opacity="0.6">
    <animate attributeName="opacity" values="0.6;1;0.6" dur="1.8s" repeatCount="indefinite"/>
  </circle>
  <circle cx="200" cy="400" r="1.1" fill="#ffffff" opacity="0.7">
    <use href="#twinkle"/>
  </circle>
  <circle cx="800" cy="450" r="1.4" fill="#ffff99" opacity="0.8">
    <animate attributeName="opacity" values="0.8;1;0.8" dur="2.2s" repeatCount="indefinite"/>
  </circle>
  <circle cx="100" cy="600" r="1" fill="#99ffcc" opacity="0.5">
    <use href="#twinkle"/>
  </circle>
  <circle cx="950" cy="650" r="1.2" fill="#ffffff" opacity="0.7">
    <animate attributeName="opacity" values="0.7;1;0.7" dur="2.8s" repeatCount="indefinite"/>
  </circle>
  
  <!-- Title -->
  <text x="561" y="80" font-family="Arial, sans-serif" font-size="48" font-weight="bold" fill="#00ffff" text-anchor="middle" filter="url(#glow)">
    COSMIC JOURNEY
  </text>
  <text x="561" y="120" font-family="Arial, sans-serif" font-size="24" fill="#ffff99" text-anchor="middle">
    ROADMAP TO THE STARS
  </text>
  
  <!-- Journey Path - CORRECTED -->
  <path d="M 150 250 Q 300 200 450 280 Q 600 350 750 300 Q 850 250 900 350 Q 950 450 800 500 Q 650 550 500 600 Q 350 650 200 750 Q 150 850 300 900 Q 450 950 600 1000 Q 750 1050 850 1150 Q 900 1250 750 1300 Q 650 1280 450 1300 Q 400 1280 350 1250 Q 300 1270 200 1300 Q 150 1350 600 1450" 
        stroke="url(#pathGrad)" 
        stroke-width="4" 
        fill="none" 
        opacity="0.8">
    <animate attributeName="stroke-dasharray" values="0,1000;1000,0" dur="8s" repeatCount="indefinite"/>
  </path>
  
  <!-- Animated Spaceship at starting point -->
  <g transform="translate(150,250)">
    <!-- Thruster glow -->
    <ellipse cx="-15" cy="0" rx="25" ry="8" fill="url(#thruster)" opacity="0.8"/>
    <!-- Spaceship body -->
    <polygon points="0,0 -20,-8 -25,-5 -25,5 -20,8 0,0 15,-3 20,0 15,3" fill="#silver" stroke="#333" stroke-width="1"/>
    <polygon points="0,0 15,-3 20,0 15,3" fill="#cccccc"/>
    <!-- Cockpit -->
    <circle cx="10" cy="0" r="4" fill="#66ccff" opacity="0.8"/>
    <!-- Animation -->
    <animateTransform attributeName="transform" type="translate" 
      values="0,0; 2,-1; 0,0; -1,1; 0,0" dur="3s" repeatCount="indefinite"/>
  </g>
  
  <!-- Planets and Destinations -->
  
  <!-- Klingon Carpark -->
  <g transform="translate(300,200)">
    <circle r="25" fill="#8B0000" filter="url(#strongGlow)"/>
    <circle r="20" fill="#DC143C"/>
    <polygon points="-8,-8 8,-8 0,8" fill="#FFD700" opacity="0.8"/>
    <text x="0" y="50" font-family="Arial, sans-serif" font-size="14" font-weight="bold" fill="#FFD700" text-anchor="middle">KLINGON</text>
    <text x="0" y="65" font-family="Arial, sans-serif" font-size="14" font-weight="bold" fill="#FFD700" text-anchor="middle">CARPARK</text>
  </g>
  
  <!-- Mount Olympus -->
  <g transform="translate(450,280)">
    <circle r="30" fill="#4169E1" filter="url(#strongGlow)"/>
    <circle r="25" fill="#6495ED"/>
    <polygon points="-10,-10 0,-20 10,-10 5,-5 -5,-5" fill="#FFFFFF" opacity="0.9"/>
    <text x="0" y="55" font-family="Arial, sans-serif" font-size="14" font-weight="bold" fill="#FFFFFF" text-anchor="middle">MOUNT</text>
    <text x="0" y="70" font-family="Arial, sans-serif" font-size="14" font-weight="bold" fill="#FFFFFF" text-anchor="middle">OLYMPUS</text>
  </g>
  
  <!-- Bowie Zone -->
  <g transform="translate(750,300)">
    <circle r="28" fill="#FF6347" filter="url(#strongGlow)"/>
    <circle r="23" fill="#FF7F50"/>
    <path d="M -15,-5 L 15,5 M -15,5 L 15,-5" stroke="#FFD700" stroke-width="3"/>
    <circle cx="0" cy="0" r="8" fill="#FFD700" opacity="0.3"/>
    <text x="0" y="50" font-family="Arial, sans-serif" font-size="14" font-weight="bold" fill="#FFD700" text-anchor="middle">BOWIE</text>
    <text x="0" y="65" font-family="Arial, sans-serif" font-size="14" font-weight="bold" fill="#FFD700" text-anchor="middle">ZONE</text>
  </g>
  
  <!-- Doge Meteor Shower -->
  <g transform="translate(900,350)">
    <circle r="26" fill="#DAA520" filter="url(#strongGlow)"/>
    <circle r="21" fill="#FFD700"/>
    <!-- Meteor streaks -->
    <line x1="-15" y1="-15" x2="-5" y2="-5" stroke="#FFFFFF" stroke-width="2" opacity="0.8">
      <animate attributeName="opacity" values="0.8;0.3;0.8" dur="1s" repeatCount="indefinite"/>
    </line>
    <line x1="8" y1="-18" x2="18" y2="-8" stroke="#FFFFFF" stroke-width="1.5" opacity="0.7">
      <animate attributeName="opacity" values="0.7;0.2;0.7" dur="1.2s" repeatCount="indefinite"/>
    </line>
    <line x1="-20" y1="5" x2="-10" y2="15" stroke="#FFFFFF" stroke-width="2" opacity="0.6">
      <animate attributeName="opacity" values="0.6;0.1;0.6" dur="0.8s" repeatCount="indefinite"/>
    </line>
    <line x1="12" y1="8" x2="22" y2="18" stroke="#FFFFFF" stroke-width="1.5" opacity="0.8">
      <animate attributeName="opacity" values="0.8;0.4;0.8" dur="1.5s" repeatCount="indefinite"/>
    </line>
    <!-- Meteor heads -->
    <circle cx="-5" cy="-5" r="2" fill="#FFFFFF" opacity="0.9">
      <animate attributeName="opacity" values="0.9;0.4;0.9" dur="1s" repeatCount="indefinite"/>
    </circle>
    <circle cx="18" cy="-8" r="1.5" fill="#FFFFFF" opacity="0.8">
      <animate attributeName="opacity" values="0.8;0.3;0.8" dur="1.2s" repeatCount="indefinite"/>
    </circle>
    <circle cx="-10" cy="15" r="2" fill="#FFFFFF" opacity="0.7">
      <animate attributeName="opacity" values="0.7;0.2;0.7" dur="0.8s" repeatCount="indefinite"/>
    </circle>
    <circle cx="22" cy="18" r="1.5" fill="#FFFFFF" opacity="0.9">
      <animate attributeName="opacity" values="0.9;0.5;0.9" dur="1.5s" repeatCount="indefinite"/>
    </circle>
    <text x="0" y="50" font-family="Arial, sans-serif" font-size="11" font-weight="bold" fill="#FFFFFF" text-anchor="middle">DOGE METEOR</text>
    <text x="0" y="65" font-family="Arial, sans-serif" font-size="11" font-weight="bold" fill="#FFFFFF" text-anchor="middle">SHOWER</text>
  </g>
  
  <!-- Planet Cyclops -->
  <g transform="translate(800,500)">
    <circle r="32" fill="#32CD32" filter="url(#strongGlow)"/>
    <circle r="27" fill="#7FFF00"/>
    <circle cx="0" cy="-5" r="12" fill="#FF0000"/>
    <circle cx="0" cy="-5" r="8" fill="#FFFFFF"/>
    <circle cx="0" cy="-5" r="4" fill="#000"/>
    <text x="0" y="55" font-family="Arial, sans-serif" font-size="14" font-weight="bold" fill="#FFFFFF" text-anchor="middle">PLANET</text>
    <text x="0" y="70" font-family="Arial, sans-serif" font-size="14" font-weight="bold" fill="#FFFFFF" text-anchor="middle">CYCLOPS</text>
  </g>
  
  <!-- Hades -->
  <g transform="translate(500,600)">
    <circle r="35" fill="#8B0000" filter="url(#strongGlow)"/>
    <circle r="30" fill="#B22222"/>
    <circle cx="-8" cy="-8" r="3" fill="#FF4500" opacity="0.8">
      <animate attributeName="r" values="3;5;3" dur="1s" repeatCount="indefinite"/>
    </circle>
    <circle cx="8" cy="-8" r="3" fill="#FF4500" opacity="0.8">
      <animate attributeName="r" values="3;5;3" dur="1.2s" repeatCount="indefinite"/>
    </circle>
    <circle cx="0" cy="8" r="4" fill="#FF4500" opacity="0.8">
      <animate attributeName="r" values="4;6;4" dur="0.8s" repeatCount="indefinite"/>
    </circle>
    <text x="0" y="60" font-family="Arial, sans-serif" font-size="16" font-weight="bold" fill="#FF4500" text-anchor="middle">HADES</text>
  </g>
  
  <!-- Planet Dad -->
  <g transform="translate(200,750)">
    <circle r="29" fill="#8B4513" filter="url(#strongGlow)"/>
    <circle r="24" fill="#D2691E"/>
    <rect x="-12" y="-15" width="24" height="8" fill="#654321" rx="2"/>
    <circle cx="-6" cy="-3" r="2" fill="#333"/>
    <circle cx="6" cy="-3" r="2" fill="#333"/>
    <rect x="-8" y="5" width="16" height="4" fill="#654321"/>
    <text x="0" y="50" font-family="Arial, sans-serif" font-size="14" font-weight="bold" fill="#FFFFFF" text-anchor="middle">PLANET</text>
    <text x="0" y="65" font-family="Arial, sans-serif" font-size="14" font-weight="bold" fill="#FFFFFF" text-anchor="middle">DAD</text>
  </g>
  
  <!-- Planet Donkey -->
  <g transform="translate(300,900)">
    <circle r="27" fill="#696969" filter="url(#strongGlow)"/>
    <circle r="22" fill="#A9A9A9"/>
    <ellipse cx="-8" cy="-10" rx="4" ry="8" fill="#654321"/>
    <ellipse cx="8" cy="-10" rx="4" ry="8" fill="#654321"/>
    <circle cx="-5" cy="0" r="2" fill="#000"/>
    <circle cx="5" cy="0" r="2" fill="#000"/>
    <ellipse cx="0" cy="8" rx="6" ry="3" fill="#FF69B4"/>
    <text x="0" y="50" font-family="Arial, sans-serif" font-size="14" font-weight="bold" fill="#FFFFFF" text-anchor="middle">PLANET</text>
    <text x="0" y="65" font-family="Arial, sans-serif" font-size="14" font-weight="bold" fill="#FFFFFF" text-anchor="middle">DONKEY</text>
  </g>
  
  <!-- Siren Solar System -->
  <g transform="translate(600,1000)">
    <circle r="20" fill="#FF1493" filter="url(#glow)"/>
    <circle r="16" fill="#FF69B4"/>
    <circle cx="25" cy="0" r="8" fill="#DA70D6" opacity="0.7">
      <animateTransform attributeName="transform" type="rotate" values="0;360" dur="4s" repeatCount="indefinite"/>
    </circle>
    <circle cx="-25" cy="0" r="6" fill="#BA55D3" opacity="0.7">
      <animateTransform attributeName="transform" type="rotate" values="360;0" dur="6s" repeatCount="indefinite"/>
    </circle>
    <path d="M -8,-4 Q 0,-8 8,-4 Q 0,0 -8,-4" fill="#FFFFFF" opacity="0.8"/>
    <text x="0" y="50" font-family="Arial, sans-serif" font-size="12" font-weight="bold" fill="#FFFFFF" text-anchor="middle">SIREN SOLAR</text>
    <text x="0" y="65" font-family="Arial, sans-serif" font-size="12" font-weight="bold" fill="#FFFFFF" text-anchor="middle">SYSTEM</text>
  </g>
  
  <!-- Deep Space -->
  <g transform="translate(850,1150)">
    <circle r="40" fill="#000000" stroke="#4B0082" stroke-width="3" filter="url(#strongGlow)"/>
    <circle r="35" fill="#191970" opacity="0.3"/>
    <circle cx="-10" cy="-10" r="2" fill="#FFFFFF" opacity="0.8">
      <animate attributeName="opacity" values="0.3;1;0.3" dur="2s" repeatCount="indefinite"/>
    </circle>
    <circle cx="12" cy="-8" r="1.5" fill="#FFFFFF" opacity="0.6">
      <animate attributeName="opacity" values="0.6;1;0.6" dur="1.5s" repeatCount="indefinite"/>
    </circle>
    <circle cx="-8" cy="10" r="1" fill="#FFFFFF" opacity="0.7">
      <animate attributeName="opacity" values="0.4;1;0.4" dur="2.5s" repeatCount="indefinite"/>
    </circle>
    <text x="0" y="65" font-family="Arial, sans-serif" font-size="16" font-weight="bold" fill="#4B0082" text-anchor="middle">DEEP</text>
    <text x="0" y="80" font-family="Arial, sans-serif" font-size="16" font-weight="bold" fill="#4B0082" text-anchor="middle">SPACE</text>
  </g>
  
  <!-- Ship of Fools -->
  <g transform="translate(750,1300)">
    <!-- Rusty spaceship hull -->
    <ellipse cx="0" cy="0" rx="30" ry="15" fill="#8B4513" stroke="#654321" stroke-width="2"/>
    <!-- Rust patches -->
    <circle cx="-15" cy="-5" r="4" fill="#A0522D" opacity="0.8"/>
    <circle cx="10" cy="8" r="3" fill="#CD853F" opacity="0.7"/>
    <circle cx="-8" cy="12" r="2" fill="#8B7355" opacity="0.6"/>
    <!-- Cockpit dome -->
    <ellipse cx="12" cy="-3" rx="8" ry="6" fill="#696969" opacity="0.6"/>
    <!-- Engine exhausts -->
    <ellipse cx="-25" cy="-6" rx="6" ry="3" fill="#444444"/>
    <ellipse cx="-25" cy="6" rx="6" ry="3" fill="#444444"/>
    <!-- Rusted details -->
    <rect x="-10" y="-2" width="20" height="4" fill="#654321" opacity="0.8"/>
    <circle cx="5" cy="-8" r="2" fill="#8B7355"/>
    <circle cx="-5" cy="10" r="1.5" fill="#A0522D"/>
    <!-- Antenna or mast -->
    <line x1="0" y1="-15" x2="0" y2="-22" stroke="#696969" stroke-width="2"/>
    <circle cx="0" cy="-22" r="2" fill="#DC143C"/>
    <text x="0" y="40" font-family="Arial, sans-serif" font-size="14" font-weight="bold" fill="#D2691E" text-anchor="middle">SHIP OF FOOLS</text>
  </g>
  
  <!-- Planet Circe -->
  <g transform="translate(450,1300)">
    <circle r="28" fill="#9932CC" filter="url(#strongGlow)"/>
    <circle r="23" fill="#BA55D3"/>
    <path d="M -12,-6 Q 0,-12 12,-6 Q 0,0 -12,-6" fill="#FFD700" opacity="0.8"/>
    <circle cx="-6" cy="6" r="2" fill="#32CD32"/>
    <circle cx="6" cy="6" r="2" fill="#FF6347"/>
    <circle cx="0" cy="12" r="2" fill="#4169E1"/>
    <text x="0" y="50" font-family="Arial, sans-serif" font-size="14" font-weight="bold" fill="#FFFFFF" text-anchor="middle">PLANET</text>
    <text x="0" y="65" font-family="Arial, sans-serif" font-size="14" font-weight="bold" fill="#FFFFFF" text-anchor="middle">CIRCE</text>
  </g>
  
  <!-- The Moon -->
  <g transform="translate(350,1250)">
    <circle r="22" fill="#C0C0C0" filter="url(#glow)"/>
    <circle r="18" fill="#E5E5E5"/>
    <circle cx="-6" cy="-4" r="3" fill="#A9A9A9" opacity="0.6"/>
    <circle cx="4" cy="-6" r="2" fill="#A9A9A9" opacity="0.6"/>
    <circle cx="-2" cy="6" r="4" fill="#A9A9A9" opacity="0.6"/>
    <circle cx="8" cy="4" r="2" fill="#A9A9A9" opacity="0.6"/>
    <text x="0" y="45" font-family="Arial, sans-serif" font-size="14" font-weight="bold" fill="#E5E5E5" text-anchor="middle">THE MOON</text>
  </g>
  
  <!-- Planet Calypso -->
  <g transform="translate(200,1300)">
    <circle r="26" fill="#008B8B" filter="url(#strongGlow)"/>
    <circle r="21" fill="#20B2AA"/>
    <path d="M -10,-8 Q 0,-12 10,-8 Q 5,-4 0,-6 Q -5,-4 -10,-8" fill="#FFFFE0" opacity="0.9"/>
    <circle cx="-5" cy="2" r="1.5" fill="#FF69B4"/>
    <circle cx="5" cy="2" r="1.5" fill="#FF69B4"/>
    <circle cx="0" cy="8" r="2" fill="#FF1493"/>
    <text x="0" y="50" font-family="Arial, sans-serif" font-size="14" font-weight="bold" fill="#FFFFFF" text-anchor="middle">PLANET</text>
    <text x="0" y="65" font-family="Arial, sans-serif" font-size="14" font-weight="bold" fill="#FFFFFF" text-anchor="middle">CALYPSO</text>
  </g>
  
  <!-- Planet Dangar (made bigger as final destination) -->
  <g transform="translate(600,1450)">
    <circle r="40" fill="#CD853F" filter="url(#strongGlow)"/>
    <circle r="35" fill="#F4A460"/>
    <rect x="-20" y="-18" width="40" height="10" fill="#8B4513" rx="5"/>
    <circle cx="-10" cy="-3" r="4" fill="#000"/>
    <circle cx="10" cy="-3" r="4" fill="#000"/>
    <rect x="-8" y="8" width="16" height="8" fill="#654321" rx="4"/>
    <polygon points="-15,20 -8,28 8,28 15,20" fill="#228B22"/>
    <!-- Crown or special marking to show it's the final destination -->
    <polygon points="-8,-25 0,-35 8,-25 4,-20 -4,-20" fill="#FFD700" opacity="0.9"/>
    <text x="0" y="65" font-family="Arial, sans-serif" font-size="16" font-weight="bold" fill="#FFFFFF" text-anchor="middle">PLANET</text>
    <text x="0" y="80" font-family="Arial, sans-serif" font-size="16" font-weight="bold" fill="#FFFFFF" text-anchor="middle">DANGAR</text>
    <text x="0" y="95" font-family="Arial, sans-serif" font-size="12" fill="#FFD700" text-anchor="middle">★ HOME ★</text>
  </g>
  
  <!-- Decorative elements -->
  <g opacity="0.3">
    <circle cx="100" cy="1000" r="60" fill="none" stroke="#4B0082" stroke-width="1" stroke-dasharray="5,5">
      <animateTransform attributeName="transform" type="rotate" values="0 100 1000;360 100 1000" dur="20s" repeatCount="indefinite"/>
    </circle>
    <circle cx="950" cy="800" r="40" fill="none" stroke="#FF6347" stroke-width="1" stroke-dasharray="3,7">
      <animateTransform attributeName="transform" type="rotate" values="360 950 800;0 950 800" dur="15s" repeatCount="indefinite"/>
    </circle>
  </g>
  
  <!-- Footer -->
  <text x="561" y="1550" font-family="Arial, sans-serif" font-size="16" fill="#00ffff" text-anchor="middle" opacity="0.8">
  </text>
</svg>